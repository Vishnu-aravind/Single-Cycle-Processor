`timescale 0.1ns/1ps
module testbench();
reg clk;
architecture arch(clk);

initial begin
    
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
    #100 clk = 0;
    #100 clk = 1;
  
  
    
    

    
end

endmodule