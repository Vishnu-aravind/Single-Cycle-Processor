module Instruction_Memory(read_addr, Instr_out);
    input [31:0]read_addr;
    output [31:0]Instr_out;
    reg [31:0]mem1[63:0];
initial begin
    mem1[0]  <= 32'b00000000000000001000001110110011; // add x7 , x1 , x0
    mem1[3]  <= 32'b00000000000001010000000010110011; // add x1 , x10 , x0
    mem1[7]  <= 32'b00000000000000111000010100110011; // add x10 , x7 , x0
    mem1[11] <= 32'b00000000000000010000001110110011; 
    mem1[15] <= 32'b00000000000001011000000100110011;
    mem1[19] <= 32'b00000000000000111000010110110011;
    mem1[23] <= 32'b00000000000000011000001110110011;
    mem1[27] <= 32'b00000000000001100000000110110011;
    mem1[31] <= 32'b00000000000000111000011000110011;
    mem1[35] <= 32'b00000000000000100000001110110011;
    mem1[39] <= 32'b00000000000001101000001000110011;
    mem1[43] <= 32'b00000000000000111000011010110011;
    mem1[47] <= 32'b00000001010000000000101100010011; //addi x22,x0,20
    mem1[51] <= 32'b01000000110110110000001110110011; //sub x7,x22,x13
    mem1[55] <= 32'b00000000001010000100010001100011; //beq x16,x17,4
    mem1[59] <= 32'b00000010100000000000101110010011; //addi x23,x0,40
    mem1[63] <= 32'b00000001100000000000110000010011; //addi x24,x0,24
 

end
assign Instr_out = mem1[read_addr];
endmodule